module twiddle_factor(
    input [7:0] i_n,
    output signed [15:0] o_real,
    output signed [15:0] o_imag
);
    logic signed [15:0]  real_value,imag_value;

    assign o_real = real_value;
    assign o_imag = imag_value;
    
    always_comb begin
        case(i_n)
           0: real_value = 16384;
1: real_value = 16379;
2: real_value = 16364;
3: real_value = 16339;
4: real_value = 16305;
5: real_value = 16260;
6: real_value = 16206;
7: real_value = 16142;
8: real_value = 16069;
9: real_value = 15985;
10: real_value = 15892;
11: real_value = 15790;
12: real_value = 15678;
13: real_value = 15557;
14: real_value = 15426;
15: real_value = 15286;
16: real_value = 15136;
17: real_value = 14978;
18: real_value = 14810;
19: real_value = 14634;
20: real_value = 14449;
21: real_value = 14255;
22: real_value = 14053;
23: real_value = 13842;
24: real_value = 13622;
25: real_value = 13395;
26: real_value = 13159;
27: real_value = 12916;
28: real_value = 12665;
29: real_value = 12406;
30: real_value = 12139;
31: real_value = 11866;
32: real_value = 11585;
33: real_value = 11297;
34: real_value = 11002;
35: real_value = 10701;
36: real_value = 10393;
37: real_value = 10079;
38: real_value = 9759;
39: real_value = 9434;
40: real_value = 9102;
41: real_value = 8765;
42: real_value = 8423;
43: real_value = 8075;
44: real_value = 7723;
45: real_value = 7366;
46: real_value = 7005;
47: real_value = 6639;
48: real_value = 6269;
49: real_value = 5896;
50: real_value = 5519;
51: real_value = 5139;
52: real_value = 4756;
53: real_value = 4369;
54: real_value = 3980;
55: real_value = 3589;
56: real_value = 3196;
57: real_value = 2801;
58: real_value = 2404;
59: real_value = 2005;
60: real_value = 1605;
61: real_value = 1205;
62: real_value = 803;
63: real_value = 402;
64: real_value = 0;
65: real_value = -402;
66: real_value = -803;
67: real_value = -1205;
68: real_value = -1605;
69: real_value = -2005;
70: real_value = -2404;
71: real_value = -2801;
72: real_value = -3196;
73: real_value = -3589;
74: real_value = -3980;
75: real_value = -4369;
76: real_value = -4756;
77: real_value = -5139;
78: real_value = -5519;
79: real_value = -5896;
80: real_value = -6269;
81: real_value = -6639;
82: real_value = -7005;
83: real_value = -7366;
84: real_value = -7723;
85: real_value = -8075;
86: real_value = -8423;
87: real_value = -8765;
88: real_value = -9102;
89: real_value = -9434;
90: real_value = -9759;
91: real_value = -10079;
92: real_value = -10393;
93: real_value = -10701;
94: real_value = -11002;
95: real_value = -11297;
96: real_value = -11585;
97: real_value = -11866;
98: real_value = -12139;
99: real_value = -12406;
100: real_value = -12665;
101: real_value = -12916;
102: real_value = -13159;
103: real_value = -13395;
104: real_value = -13622;
105: real_value = -13842;
106: real_value = -14053;
107: real_value = -14255;
108: real_value = -14449;
109: real_value = -14634;
110: real_value = -14810;
111: real_value = -14978;
112: real_value = -15136;
113: real_value = -15286;
114: real_value = -15426;
115: real_value = -15557;
116: real_value = -15678;
117: real_value = -15790;
118: real_value = -15892;
119: real_value = -15985;
120: real_value = -16069;
121: real_value = -16142;
122: real_value = -16206;
123: real_value = -16260;
124: real_value = -16305;
125: real_value = -16339;
126: real_value = -16364;
127: real_value = -16379;
128: real_value = -16384;
129: real_value = -16379;
130: real_value = -16364;
131: real_value = -16339;
132: real_value = -16305;
133: real_value = -16260;
134: real_value = -16206;
135: real_value = -16142;
136: real_value = -16069;
137: real_value = -15985;
138: real_value = -15892;
139: real_value = -15790;
140: real_value = -15678;
141: real_value = -15557;
142: real_value = -15426;
143: real_value = -15286;
144: real_value = -15136;
145: real_value = -14978;
146: real_value = -14810;
147: real_value = -14634;
148: real_value = -14449;
149: real_value = -14255;
150: real_value = -14053;
151: real_value = -13842;
152: real_value = -13622;
153: real_value = -13395;
154: real_value = -13159;
155: real_value = -12916;
156: real_value = -12665;
157: real_value = -12406;
158: real_value = -12139;
159: real_value = -11866;
160: real_value = -11585;
161: real_value = -11297;
162: real_value = -11002;
163: real_value = -10701;
164: real_value = -10393;
165: real_value = -10079;
166: real_value = -9759;
167: real_value = -9434;
168: real_value = -9102;
169: real_value = -8765;
170: real_value = -8423;
171: real_value = -8075;
172: real_value = -7723;
173: real_value = -7366;
174: real_value = -7005;
175: real_value = -6639;
176: real_value = -6269;
177: real_value = -5896;
178: real_value = -5519;
179: real_value = -5139;
180: real_value = -4756;
181: real_value = -4369;
182: real_value = -3980;
183: real_value = -3589;
184: real_value = -3196;
185: real_value = -2801;
186: real_value = -2404;
187: real_value = -2005;
188: real_value = -1605;
189: real_value = -1205;
190: real_value = -803;
191: real_value = -402;
192: real_value = 0;
193: real_value = 402;
194: real_value = 803;
195: real_value = 1205;
196: real_value = 1605;
197: real_value = 2005;
198: real_value = 2404;
199: real_value = 2801;
200: real_value = 3196;
201: real_value = 3589;
202: real_value = 3980;
203: real_value = 4369;
204: real_value = 4756;
205: real_value = 5139;
206: real_value = 5519;
207: real_value = 5896;
208: real_value = 6269;
209: real_value = 6639;
210: real_value = 7005;
211: real_value = 7366;
212: real_value = 7723;
213: real_value = 8075;
214: real_value = 8423;
215: real_value = 8765;
216: real_value = 9102;
217: real_value = 9434;
218: real_value = 9759;
219: real_value = 10079;
220: real_value = 10393;
221: real_value = 10701;
222: real_value = 11002;
223: real_value = 11297;
224: real_value = 11585;
225: real_value = 11866;
226: real_value = 12139;
227: real_value = 12406;
228: real_value = 12665;
229: real_value = 12916;
230: real_value = 13159;
231: real_value = 13395;
232: real_value = 13622;
233: real_value = 13842;
234: real_value = 14053;
235: real_value = 14255;
236: real_value = 14449;
237: real_value = 14634;
238: real_value = 14810;
239: real_value = 14978;
240: real_value = 15136;
241: real_value = 15286;
242: real_value = 15426;
243: real_value = 15557;
244: real_value = 15678;
245: real_value = 15790;
246: real_value = 15892;
247: real_value = 15985;
248: real_value = 16069;
249: real_value = 16142;
250: real_value = 16206;
251: real_value = 16260;
252: real_value = 16305;
253: real_value = 16339;
254: real_value = 16364;
255: real_value = 16379;
            default: real_value = 0;
        endcase
    end
    always_comb begin
        case(i_n)
            0: imag_value = 0;
1: imag_value = -402;
2: imag_value = -803;
3: imag_value = -1205;
4: imag_value = -1605;
5: imag_value = -2005;
6: imag_value = -2404;
7: imag_value = -2801;
8: imag_value = -3196;
9: imag_value = -3589;
10: imag_value = -3980;
11: imag_value = -4369;
12: imag_value = -4756;
13: imag_value = -5139;
14: imag_value = -5519;
15: imag_value = -5896;
16: imag_value = -6269;
17: imag_value = -6639;
18: imag_value = -7005;
19: imag_value = -7366;
20: imag_value = -7723;
21: imag_value = -8075;
22: imag_value = -8423;
23: imag_value = -8765;
24: imag_value = -9102;
25: imag_value = -9434;
26: imag_value = -9759;
27: imag_value = -10079;
28: imag_value = -10393;
29: imag_value = -10701;
30: imag_value = -11002;
31: imag_value = -11297;
32: imag_value = -11585;
33: imag_value = -11866;
34: imag_value = -12139;
35: imag_value = -12406;
36: imag_value = -12665;
37: imag_value = -12916;
38: imag_value = -13159;
39: imag_value = -13395;
40: imag_value = -13622;
41: imag_value = -13842;
42: imag_value = -14053;
43: imag_value = -14255;
44: imag_value = -14449;
45: imag_value = -14634;
46: imag_value = -14810;
47: imag_value = -14978;
48: imag_value = -15136;
49: imag_value = -15286;
50: imag_value = -15426;
51: imag_value = -15557;
52: imag_value = -15678;
53: imag_value = -15790;
54: imag_value = -15892;
55: imag_value = -15985;
56: imag_value = -16069;
57: imag_value = -16142;
58: imag_value = -16206;
59: imag_value = -16260;
60: imag_value = -16305;
61: imag_value = -16339;
62: imag_value = -16364;
63: imag_value = -16379;
64: imag_value = -16384;
65: imag_value = -16379;
66: imag_value = -16364;
67: imag_value = -16339;
68: imag_value = -16305;
69: imag_value = -16260;
70: imag_value = -16206;
71: imag_value = -16142;
72: imag_value = -16069;
73: imag_value = -15985;
74: imag_value = -15892;
75: imag_value = -15790;
76: imag_value = -15678;
77: imag_value = -15557;
78: imag_value = -15426;
79: imag_value = -15286;
80: imag_value = -15136;
81: imag_value = -14978;
82: imag_value = -14810;
83: imag_value = -14634;
84: imag_value = -14449;
85: imag_value = -14255;
86: imag_value = -14053;
87: imag_value = -13842;
88: imag_value = -13622;
89: imag_value = -13395;
90: imag_value = -13159;
91: imag_value = -12916;
92: imag_value = -12665;
93: imag_value = -12406;
94: imag_value = -12139;
95: imag_value = -11866;
96: imag_value = -11585;
97: imag_value = -11297;
98: imag_value = -11002;
99: imag_value = -10701;
100: imag_value = -10393;
101: imag_value = -10079;
102: imag_value = -9759;
103: imag_value = -9434;
104: imag_value = -9102;
105: imag_value = -8765;
106: imag_value = -8423;
107: imag_value = -8075;
108: imag_value = -7723;
109: imag_value = -7366;
110: imag_value = -7005;
111: imag_value = -6639;
112: imag_value = -6269;
113: imag_value = -5896;
114: imag_value = -5519;
115: imag_value = -5139;
116: imag_value = -4756;
117: imag_value = -4369;
118: imag_value = -3980;
119: imag_value = -3589;
120: imag_value = -3196;
121: imag_value = -2801;
122: imag_value = -2404;
123: imag_value = -2005;
124: imag_value = -1605;
125: imag_value = -1205;
126: imag_value = -803;
127: imag_value = -402;
128: imag_value = 0;
129: imag_value = 402;
130: imag_value = 803;
131: imag_value = 1205;
132: imag_value = 1605;
133: imag_value = 2005;
134: imag_value = 2404;
135: imag_value = 2801;
136: imag_value = 3196;
137: imag_value = 3589;
138: imag_value = 3980;
139: imag_value = 4369;
140: imag_value = 4756;
141: imag_value = 5139;
142: imag_value = 5519;
143: imag_value = 5896;
144: imag_value = 6269;
145: imag_value = 6639;
146: imag_value = 7005;
147: imag_value = 7366;
148: imag_value = 7723;
149: imag_value = 8075;
150: imag_value = 8423;
151: imag_value = 8765;
152: imag_value = 9102;
153: imag_value = 9434;
154: imag_value = 9759;
155: imag_value = 10079;
156: imag_value = 10393;
157: imag_value = 10701;
158: imag_value = 11002;
159: imag_value = 11297;
160: imag_value = 11585;
161: imag_value = 11866;
162: imag_value = 12139;
163: imag_value = 12406;
164: imag_value = 12665;
165: imag_value = 12916;
166: imag_value = 13159;
167: imag_value = 13395;
168: imag_value = 13622;
169: imag_value = 13842;
170: imag_value = 14053;
171: imag_value = 14255;
172: imag_value = 14449;
173: imag_value = 14634;
174: imag_value = 14810;
175: imag_value = 14978;
176: imag_value = 15136;
177: imag_value = 15286;
178: imag_value = 15426;
179: imag_value = 15557;
180: imag_value = 15678;
181: imag_value = 15790;
182: imag_value = 15892;
183: imag_value = 15985;
184: imag_value = 16069;
185: imag_value = 16142;
186: imag_value = 16206;
187: imag_value = 16260;
188: imag_value = 16305;
189: imag_value = 16339;
190: imag_value = 16364;
191: imag_value = 16379;
192: imag_value = 16384;
193: imag_value = 16379;
194: imag_value = 16364;
195: imag_value = 16339;
196: imag_value = 16305;
197: imag_value = 16260;
198: imag_value = 16206;
199: imag_value = 16142;
200: imag_value = 16069;
201: imag_value = 15985;
202: imag_value = 15892;
203: imag_value = 15790;
204: imag_value = 15678;
205: imag_value = 15557;
206: imag_value = 15426;
207: imag_value = 15286;
208: imag_value = 15136;
209: imag_value = 14978;
210: imag_value = 14810;
211: imag_value = 14634;
212: imag_value = 14449;
213: imag_value = 14255;
214: imag_value = 14053;
215: imag_value = 13842;
216: imag_value = 13622;
217: imag_value = 13395;
218: imag_value = 13159;
219: imag_value = 12916;
220: imag_value = 12665;
221: imag_value = 12406;
222: imag_value = 12139;
223: imag_value = 11866;
224: imag_value = 11585;
225: imag_value = 11297;
226: imag_value = 11002;
227: imag_value = 10701;
228: imag_value = 10393;
229: imag_value = 10079;
230: imag_value = 9759;
231: imag_value = 9434;
232: imag_value = 9102;
233: imag_value = 8765;
234: imag_value = 8423;
235: imag_value = 8075;
236: imag_value = 7723;
237: imag_value = 7366;
238: imag_value = 7005;
239: imag_value = 6639;
240: imag_value = 6269;
241: imag_value = 5896;
242: imag_value = 5519;
243: imag_value = 5139;
244: imag_value = 4756;
245: imag_value = 4369;
246: imag_value = 3980;
247: imag_value = 3589;
248: imag_value = 3196;
249: imag_value = 2801;
250: imag_value = 2404;
251: imag_value = 2005;
252: imag_value = 1605;
253: imag_value = 1205;
254: imag_value = 803;
255: imag_value = 402;
            default: imag_value = 0;
        endcase 
    end
endmodule
